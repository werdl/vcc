module main

fn main() {
	println(lex("int main() { return 3 }"))
}
